module CPU( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset // @[:@30.4]
);
  initial begin end
endmodule
