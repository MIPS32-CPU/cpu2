module MEM( // @[:@3.2]
  input   clock, // @[:@4.4]
  input   reset // @[:@5.4]
);
  initial begin end
endmodule
